`timescale 1ns/1ns

module ROM (addr,data);
input [31:0] addr;
output [31:0] data;
reg [31:0] data;
localparam ROM_SIZE = 32;
reg [31:0] ROM_DATA[ROM_SIZE-1:0];

always@(*)
	case(addr[9:2])	//Address Must Be Word Aligned.
0:	data <= 32'b00001000000000000000000000000011;
1:	data <= 32'b00001000000000000000000000110001;
2:	data <= 32'b00001000000000000000000010001111;
3:	data <= 32'b00000000000000001110100000100000;
4:	data <= 32'b00111100000101110100000000000000;
5:	data <= 32'b00000000000000001011000000100111;
6:	data <= 32'b10101110111000000000000000001100;
7:	data <= 32'b10101110111101100000000000010100;
8:	data <= 32'b10101110111000000000000000001000;
9:	data <= 32'b00100010110010001001111001011000;
10:	data <= 32'b00100001000010001001111001011000;
11:	data <= 32'b10101110111010000000000000000000;
12:	data <= 32'b10101110111101100000000000000100;
13:	data <= 32'b00100000000010000000000000000011;
14:	data <= 32'b10101110111010000000000000001000;
15:	data <= 32'b10101110111010000000000000100000;
16:	data <= 32'b00000000000000001000000000100000;
17:	data <= 32'b00000000000000000000000000000000;
18:	data <= 32'b10001110111010000000000000100000;
19:	data <= 32'b00100000000010010000000000001000;
20:	data <= 32'b00000001001010000101000000100100;
21:	data <= 32'b00010001010000001111111111111100;
22:	data <= 32'b00010110000000000000000000000011;
23:	data <= 32'b10001110111001000000000000011100;
24:	data <= 32'b00100000000100000000000000000001;
25:	data <= 32'b00001000000000000000000000010010;
26:	data <= 32'b10001110111001010000000000011100;
27:	data <= 32'b00001100000000000000000000100101;
28:	data <= 32'b00000000000000001000000000100000;
29:	data <= 32'b10101110111000100000000000001100;
30:	data <= 32'b10001110111010000000000000100000;
31:	data <= 32'b00100000000010010000000000010000;
32:	data <= 32'b00000001000010010101000000100100;
33:	data <= 32'b00000000000010100101000100000010;
34:	data <= 32'b00010101010000001111111111111011;
35:	data <= 32'b10101110111000100000000000011000;
36:	data <= 32'b00001000000000000000000000010010;
37:	data <= 32'b00000000100000000100000000100000;
38:	data <= 32'b00000000101000000100100000100000;
39:	data <= 32'b00010001000010010000000000000111;
40:	data <= 32'b00000001000010010101000000100010;
41:	data <= 32'b00011101010000000000000000000011;
42:	data <= 32'b00000001000000000101000000100000;
43:	data <= 32'b00000001001000000100000000100000;
44:	data <= 32'b00000001010000000100100000100000;
45:	data <= 32'b00000001000010010100000000100010;
46:	data <= 32'b00001000000000000000000000100111;
47:	data <= 32'b00000001000000000001000000100000;
48:	data <= 32'b00000011111000000000000000001000;
49:	data <= 32'b10001110111101010000000000001000;
50:	data <= 32'b00100010110101001111111111111010;
51:	data <= 32'b00000010100101011010100000100100;
52:	data <= 32'b10101110111101010000000000001000;
53:	data <= 32'b10101111101010000000000000000000;
54:	data <= 32'b10101111101010010000000000000100;
55:	data <= 32'b10101111101010100000000000001000;
56:	data <= 32'b10101111101010110000000000001100;
57:	data <= 32'b10101111101011000000000000010000;
58:	data <= 32'b10101111101011010000000000010100;
59:	data <= 32'b00100011101111010000000000010100;
60:	data <= 32'b10001110111010000000000000010100;
61:	data <= 32'b00000000000010000100001000000010;
62:	data <= 32'b00110000100010010000000011110000;
63:	data <= 32'b00000000000010010100100100000010;
64:	data <= 32'b00100000000010100000000000001110;
65:	data <= 32'b00100000000010110000000000000111;
66:	data <= 32'b00010001000010100000000000001101;
67:	data <= 32'b00110000100010010000000000001111;
68:	data <= 32'b00100000000010100000000000000111;
69:	data <= 32'b00100000000010110000000000001011;
70:	data <= 32'b00010001000010100000000000001001;
71:	data <= 32'b00110000101010010000000011110000;
72:	data <= 32'b00000000000010010100100100000010;
73:	data <= 32'b00100000000010100000000000001011;
74:	data <= 32'b00100000000010110000000000001101;
75:	data <= 32'b00010001000010100000000000000100;
76:	data <= 32'b00110000101010010000000000001111;
77:	data <= 32'b00100000000010100000000000001101;
78:	data <= 32'b00100000000010110000000000001110;
79:	data <= 32'b00010001000010100000000000000000;
80:	data <= 32'b00100000000011000000000011000000;
81:	data <= 32'b00100000000011010000000000000000;
82:	data <= 32'b00010001001011010000000000101101;
83:	data <= 32'b00100000000011000000000011111001;
84:	data <= 32'b00100000000011010000000000000001;
85:	data <= 32'b00010001001011010000000000101010;
86:	data <= 32'b00100000000011000000000010100100;
87:	data <= 32'b00100000000011010000000000000010;
88:	data <= 32'b00010001001011010000000000100111;
89:	data <= 32'b00100000000011000000000010110000;
90:	data <= 32'b00100000000011010000000000000011;
91:	data <= 32'b00010001001011010000000000100100;
92:	data <= 32'b00100000000011000000000010011001;
93:	data <= 32'b00100000000011010000000000000100;
94:	data <= 32'b00010001001011010000000000100001;
95:	data <= 32'b00100000000011000000000010010010;
96:	data <= 32'b00100000000011010000000000000101;
97:	data <= 32'b00010001001011010000000000011110;
98:	data <= 32'b00100000000011000000000010000010;
99:	data <= 32'b00100000000011010000000000000110;
100:	data <= 32'b00010001001011010000000000011011;
101:	data <= 32'b00100000000011000000000011111000;
102:	data <= 32'b00100000000011010000000000000111;
103:	data <= 32'b00010001001011010000000000011000;
104:	data <= 32'b00100000000011000000000010000000;
105:	data <= 32'b00100000000011010000000000001000;
106:	data <= 32'b00010001001011010000000000010101;
107:	data <= 32'b00100000000011000000000010010000;
108:	data <= 32'b00100000000011010000000000001001;
109:	data <= 32'b00010001001011010000000000010010;
110:	data <= 32'b00100000000011000000000010001000;
111:	data <= 32'b00100000000011010000000000001010;
112:	data <= 32'b00010001001011010000000000001111;
113:	data <= 32'b00100000000011000000000010000011;
114:	data <= 32'b00100000000011010000000000001011;
115:	data <= 32'b00010001001011010000000000001100;
116:	data <= 32'b00100000000011000000000011000110;
117:	data <= 32'b00100000000011010000000000001100;
118:	data <= 32'b00010001001011010000000000001001;
119:	data <= 32'b00100000000011000000000010100001;
120:	data <= 32'b00100000000011010000000000001101;
121:	data <= 32'b00010001001011010000000000000110;
122:	data <= 32'b00100000000011000000000010000110;
123:	data <= 32'b00100000000011010000000000001110;
124:	data <= 32'b00010001001011010000000000000011;
125:	data <= 32'b00100000000011000000000010001110;
126:	data <= 32'b00100000000011010000000000001111;
127:	data <= 32'b00010001001011010000000000000000;
128:	data <= 32'b00000000000010110101101000000000;
129:	data <= 32'b00000001011011000100000000100000;
130:	data <= 32'b10101110111010000000000000010100;
131:	data <= 32'b10001111101011010000000000000000;
132:	data <= 32'b10001111101011001111111111111100;
133:	data <= 32'b10001111101010111111111111111000;
134:	data <= 32'b10001111101010101111111111110100;
135:	data <= 32'b10001111101010011111111111110000;
136:	data <= 32'b10001111101010001111111111101100;
137:	data <= 32'b00100011101111011111111111101100;
138:	data <= 32'b10001110111101010000000000001000;
139:	data <= 32'b00100000000101000000000000000010;
140:	data <= 32'b00000010100101011010100000100101;
141:	data <= 32'b10101110111101010000000000001000;
142:	data <= 32'b00000011010000000000000000001000;
143:	data <= 32'b00000000000000000000000000000000;


	   default:	data <= 32'b00000011010000000000000000001000;
	endcase
endmodule
